work.mem(main) :8: :4:
